* D:\LTspiceWorldTour2009\4884.asc
XX1 N001 N002 0 SI4884DY
V1 N001 0 0
V2 N002 0 0
.dc V1 0 10 2m V2 4 8 2
*$
.SUBCKT SI4884DY 4 1 2
M1  3 1 2 2 NMOS W=3185952u L=0.50u 
M2  2 1 2 4 PMOS W=3185952u L=0.34u
R1  4 3     RTEMP 49E-4
CGS 1 2     720E-12
DBD 2 4     DBD
**************************************************************************************************
.MODEL NMOS NMOS(LEVEL = 3    TOX  = 5E-8    RS    = 22E-4 NSUB  = 17E16
+ KP   = 1.3E-5  UO   = 650   VMAX = 0       XJ    = 5E-7  KAPPA = 25E-2
+ ETA  = 1E-4    TPG  = 1     IS   = 0       LD    = 0     CGSO  = 0
+ CGDO = 0       CGBO = 0     NFS  = 0.8E12  DELTA = 0.1)
*************************************************************************************************
.MODEL PMOS PMOS(LEVEL = 3  TOX = 5E-8   NSUB = 1.95E16   TPG = -1) 
*************************************************************************************************
.MODEL DBD D(CJO=1.1n VJ=.38 M=.32 RS=.035 FC=.5 IS=1E-11 TT=30n N=1 BV=50)
*************************************************************************************************
.MODEL RTEMP RES(TC1=6.5E-3 TC2=5.5E-6)
*************************************************************************************************
.ENDS
.probe
.end
