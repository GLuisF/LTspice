DGMOSTST
**********
.OP
.INCLUDE DG_MOS.LIB
*MAKE SURE TO USE THE CORRECT .LIB FILENAME 
*DEFINE DUT=MN201
*REPLACE DUT= WITH DUT=YOUR MODEL NAME
*FOR P CHANNEL FETS FLIP VGS, VDS, AND V2
.DC VDS 0 20 .1 VGS1 -1 1 .5 
*.DC VGS1 -1.5 1 .1 VGS2 0 4 1 
*FOR ID VS. VGS CURVE, USE .DC VGS ONLY, PLOT I(V3) VS. VGS
*SPICE_NET
*ALIAS  I(V3)=ID
.PRINT DC  I(V3)
VDS 4 0 15
*SET VDS RANGE IN THE .DC STATEMENT 
VGS2 1 0 4
*SET VGS RANGE IN THE .DC STATEMENT 
X3 5 1 3 0 MN201
V6 3 2 
VGS1 2 0 
V3 4 5 
.END
