* This subcircuit models an opamp in a circuit
* OPamp Inverting circuit
 
* subcirciut of internal connections of opamp
.SUBCKT Opamp p_in n_in com out
EX int com p_in n_in 1e5
Ri p_in n_in 500K
Ro int out 50.0
.ENDS
 
* circuit elements connected to opamp
 
Vg 1 0 DC 50mV
Rg 1 2 5K
Rf 2 3 50K
Rl 3 0 20K
X1 0 2 0 3 opamp

.OP 
*.DC Vg 50m 50m 1m ; No sweep only one point
.END
