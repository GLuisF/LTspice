*
L1 N001 0 Flux=tanh(x) ; x is a keyword for the current
I1 0 N001 PWL(0 0 10 10)
.tran 5
.end
