* AD746 SPICE Macro-model       		3/91, Rev. B
*                                               JLW / PMI
*
* Revision History:
*     Corrected VOS to be 0.25mV
*
*
* This version of the AD746 model simulates the typical
* parameters corresponding to those in the device data
* sheet.
*
*
* Copyright 1991 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* connections: non-inverting input
*               |  inverting input
*               |  |  positive power supply
*               |  |  |  negative power supply
*               |  |  |  |  output
*               |  |  |  |  | 
.subckt AD746  11 14 10 16 13 
* 
VOS 14 7 DC 0.25E-3
EC 8 0 (13,0) 1
C1 5 6 0.33E-12
GB 12 0 (15,0) 1.67E3 
RD1 5 16 16E3
RD2 6 16 16E3
ISS 10 1 DC 100E-6
GCM 0 15 (0,1) 1.76E-9
GA 15 0 (6,5) 1.75E-3
RE 1 0 2.5E6
RGM 15 0 1.76E3
VC 10 2 DC 2.8
VE 9 16 DC 2.8
RO1 12 13 25
CE 1 0 1E-12
RO2 0 12 30
RS1 1 3 5.77E3
RS2 1 4 5.77E3
CCI 15 12 40E-12
RP 16 10 8.5E3
J1 5 11 3 FET
J2 6 7 4 FET
DC 13 2 DIODE
DE 9 13 DIODE
DP 16 10 DIODE
D1 8 12 DIODE
D2 12 8 DIODE
.MODEL DIODE D()
.MODEL FET PJF(VTO=-1 BETA=1E-3 IS=110E-12)
.ENDS
