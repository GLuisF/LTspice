* d:\Arrow\astable.asc
R1 N001 N002 2K
R2 N001 N003 2K
R3 N002 N004 101K
R4 N003 N005 100K
C1 N003 N004 .01�
C2 N005 N002 .01�
V1 N001 0 5
Q1 N003 N005 0 0 2N3904
Q2 N002 N004 0 0 2N3904
.lib C:\LTspice\lib\cmp\standard.bjt
.tran 25m startup
.end
