* C:\Archivos de programa\LTC\SwCADIII\examples\Robertugo\Convert\Tero\Tero555ALL.asc
Ct N001 0 820p
DretInv 0 N003 1N914
Dalim Out Alim555 MURS120
Dpol N005 N004 MBRS1100
Rtoff N001 N002 47K tol=1 pwr=0.1
Rton Alim555 N002 27K tol=1 pwr=0.1
QCtrl PwmCtrl beQctrl 0 0 BC547A
Rd2 beQctrl 0 1K tol=1 pwr=0.1
VLocom N006 0 80v AC 1 Rser=1m
RDis N004 Alim555 22k tol=10 pwr=5
R_uFan Alim555 0 150 tol=1 pwr=0.1
Rbuf N003 Out_555 47 tol=1 pwr=0.1
Rbmin N003 0 22 tol=1 pwr=0.1
Cf1 OutRect 0 220� V=16 Irms=2.4 Rser=0.05 MTBF=0 Lser=2.1p ppPkg=1
Cf2 Out 0 220� V=16 Irms=2.4 Rser=0.05 MTBF=0 Lser=2.1p ppPkg=1
Lf Out OutRect 100� Ipk=10 Rser=0.001 Rpar=0 Cpar=0
Cstart N004 Alim555 47� V=100 Irms=210m Rser=0.37 MTBF=2000 Lser=0 mfg="Nichicon" pn="UPR2A470MPH" type="Al electrolytic" ppPkg=1
Csnub High 0 1n2 Rser=10
D2 N002 N001 1N914
LP N004 High 904� Rser=1 Rpar=1430 Cpar=5p
LS 0 N007 50� Rser=0.01 Rpar=110
Drect N007 OutRect MBR735
Qout High N003 0 0 BU508
XU1 0 N001 Out_555 Alim555 PwmCtrl N001 N002 Alim555 NE555
Csint N007 0 {100n}
Rd1 beQctrl OutRect 18K tol=1 pwr=0.1
Rlim N005 N006 2R2 tol=1 pwr=0.1
Cps N007 High 10p
Cf3 Alim555 0 220� V=16 Irms=2.4 Rser=0.05 MTBF=0 Lser=2.1p ppPkg=1
iLoad Out 0 3
.model D D
.lib 'C:\Archivos de programa\LTC\SwCADIII\lib\cmp\standard.dio'
.model NPN NPN
.model PNP PNP
.lib 'C:\Archivos de programa\LTC\SwCADIII\lib\cmp\standard.bjt'
K1 LP LS .995
.tran 0 5m startup
* (18K)
* x100V
* x250V
* 2R7min
* Varilla de ferrite,\nbobinada a tope.\nLargo=50mm,\ndi�metro=8mm.\nLP=904uH=170esp,\ndiam=0.25mm.\nLS=50uH=40esp. y\ndiam=1mm.
* Cheap & dirty(some\nfreq var) for 80V\n(Locomotive) to\n12V x 3A PWM\n  Flyback. If short-\n  circuit autostop!\n  Ef(35W)>70%\n  &Full NE555\n  bipolar use.
* El modelo TLC555 de Helmut, no funciona correctamente; (problemas con Ctrl).
* .step param val 80n 120n 20n
* 56K
* 22K
.lib 'C:\Archivos de programa\LTC\SwCADIII\lib\sub\timers.lib'
.backanno
.end
