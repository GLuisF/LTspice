* Verilog-A vbic_3T_it_cf test circuit
vbe bx 0 0
vcb cx bx 0
vib bx b 0
vic cx c 0
q1 c b 0 vbic
.model vbic npn(level=9 RCX=10 RCI=10 RBX=1 RBI=10 RE=1 RBP=10 RS=10
IBEN=1.0e-13 RTH=100)
.dc vbe 0.5 1.0 0.001
.probe i(vib) i(vic)
.end