* AD626 SPICE Macro-model               Rev. A, 11/95
*                                       ARG / ADSC
*
* Copyright 1995 by Analog Devices
*
* Refer to "README.DOC" file for License Statement. Use of
* this model indicates your acceptance of the terms and pro-
* visions in the License Statement.
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  gain=100
*                |  |  |  |  |  filter
*                |  |  |  |  |  |  ground
*                |  |  |  |  |  |  |  output
*                |  |  |  |  |  |  |  |
.SUBCKT AD626    1  2  99 50 30 31 90 49
*
* A1 INPUT ATTENUATORS, GAIN, AND OFFSET RESISTORS
*
R1 1 3 200K
R2 2 4 200K
RS1 3 16 1K
RS2 4 18 1K
R3 3 5 41K
R4 4 6 41K
R5 5 6 4.244K TC=-13.4U
R6 5 0 540
R7 6 0 540
R9 6 7 10K
R11 5 0 10K
C1 16 0 5P
C2 17 0 5P
*
* A1 INPUT STAGE AND POLE AT 1MHZ
*
I1 99 8 7.55U
Q1 11 16 9 QP 1
Q2 12 17 10 QP 1
R21 11 50 13.7934K
R22 12 50 13.7934K
R23 8 9 6.89705K
R24 8 10 6.89705K
C3 11 12 5.769P
EOS 61 17 POLY(1) 33 98 1.43U 0.537
ETC 18 61 POLY(1) 60 0 -49.665M 1
ITC 0 60 49.665U
RTC 60 0 1K TC=-81.8U
*
* GAIN STAGE AND DOMINANT POLE AT 120HZ
*
EREF 98 0 POLY(2) 99 0 50 0 0 0.5 0.5
G1 98 13 12 11 72.4983U
R25 13 98 13.7934E6
C4 13 98 96.154P
D1 13 99 DX
D2 50 13 DX
*
* COMMON MODE STAGE WITH ZERO AT 1.78KHZ
*
ECM 32 98 POLY(2) 1 98 2 98 0 0.5 0.5
R28 32 33 1E6
R29 33 98 10
CCM 32 33 503P
*
* NEGATIVE ZERO AT 0.6MHZ
*
E1 23 98 13 98 1E6
R26 23 24 1E3
R27 24 98 1E-3
FNZ 23 24 VNZ -1
ENZ 25 98 23 24 1
VNZ 26 98 DC 0
CNZ 25 26 265P
*
* POLE AT 5MHZ
*
G2 98 20 24 98 1E-6
R30 20 98 1E6
C5 20 98 32F
*
* A1 OUTPUT STAGE
*
EIN1 99 27 POLY(1) 20 98 1.5102 1.124
Q216 50 27 28 QP375 3.444
Q218 7 29 99 QP350 9.913
R31 28 29 27K
I2 99 29 4.75U
R8 7 50 10K
R12 7 31 100K
*
* A2 INPUT STAGE
*
I3 99 34 2.516667U
Q3 35 31 37 QP 1
Q4 36 39 38 QP 1
R32 35 50 106.103K
R33 36 50 106.103K
R34 34 37 85.414K
R35 34 38 85.414K
R10 41 0 10K
R13 49 50 10K
R14 41 30 555.71 TC=-4.5U
R15 41 49 10K
R17 39 41 95K
*
* A2 1ST GAIN STAGE AND SLEW RATE
*
G3 98 42 36 35 30.159U
R36 42 98 1E6
E2 99 43 POLY(1) 99 98 -0.473 1
E3 44 50 POLY(1) 98 50 -0.473 1
D3 42 43 DX
D4 44 42 DX
*
* A2 2ND GAIN STAGE AND DOMINANT POLE AT 12HZ
*
G4 98 45 42 98 2.5U
R37 45 98 132.629E6
C7 45 98 100P
D5 45 59 DX
D6 55 45 DX
VC1 59 99 5
VC2 50 55 5
*
* NEGATIVE ZERO AT 1MHZ
*
E4 51 98 45 98 1E6
R38 51 52 1E6
R39 52 98 1
FNZ2 51 52 VNZ2 -1
ENZ2 53 98 51 52 1
VNZ2 54 98 0
CNZ2 53 54 159F
*
* A2 OUTPUT STAGE
*
GSY 99 50 99 50 29.2U
EIN2 99 56 POLY(1) 52 98 1.75608 46.605E-3
RIN 46 56 10K
Q316 50 46 47 QP375 1.778
Q310 50 47 48 QP375 5.925
Q318 49 48 57 50 QP350 9.913
I4 99 47 4.75U
I5 99 48 9.5U
VSC 99 57 0.03
FSC 58 99 VSC 1
QSC 46 58 99 QP350 1
RSC 99 58 48
*
* MODELS USED
*
.MODEL QP350 PNP(IS=1.4E-15 BF=70 CJE=.012P CJC=.06P RE=20 RB=350
+RC=200)
.MODEL QP375 PNP(IS=1.4E-15 CJE=.01P CJC=.05P RE=20 RC=400 RB=100)
.MODEL QP AKO:QP350 PNP(BF=150 VA=100)
.MODEL DX D(CJO=1F RS=.1)
.ENDS
