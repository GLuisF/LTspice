.SUBCKT irf7343 1 2 3 4 6 8
* DUAL N AND P CHANNEL MOSFET
* External Node Designations
* Node 1 -> N-channel Source
* Node 2 -> N-Channel Gate
* Node 3 -> P-Channel Source
* Node 4 -> P-Channel Gate
* Node 6 -> P-Channel Drain
* Node 8 -> N-Channel Drain
X1 8 2 1 irf7343-n-ch
X2 6 4 3 irf7343-p-ch
.ENDS irf7343

.SUBCKT irf7343-n-ch 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Mar 22, 04
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=2.21828 LAMBDA=0 KP=31.0598
+CGSO=6.94399e-06 CGDO=4.54721e-07
RS 8 3 0.0239533
D1 3 1 MD
.MODEL MD D IS=4.51343e-09 RS=0.00912834 N=1.5 BV=55
+IBV=0.00025 EG=1.2 XTI=2.93898 TT=1.0e-07
+CJO=5.06742e-10 VJ=1.604 M=0.497938 FC=0.5
RDS 3 1 1e+06
RD 9 1 0.0177251
RG 2 7 1.70427
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=8.4332e-10 VJ=0.500018 M=0.882099 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.408289 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 1.15932e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.408289
.ENDS irf7343-n-ch

.SUBCKT irf7343-p-ch 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Mar 23, 04
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM PMOS LEVEL=1 IS=1e-32
+VTO=-2.19655 LAMBDA=0.00706611 KP=6.18356
+CGSO=6.43304e-06 CGDO=4.93008e-07
RS 8 3 0.0484461
D1 1 3 MD
.MODEL MD D IS=1.58336e-10 RS=0.0175907 N=1.27607 BV=55
+IBV=0.00025 EG=1 XTI=4 TT=-1.0e-07
+CJO=6.06157e-10 VJ=0.812982 M=0.454501 FC=0.1
RDS 3 1 1e+06
RD 9 1 0.0292188
RG 2 7 6.30602
D2 5 4 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=8.92291e-10 VJ=0.5 M=0.817556 FC=1e-08
D3 5 0 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.400161 RS=3.00001e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 1.35866e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 6 0 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.400161
.ENDS irf7343-p-ch

