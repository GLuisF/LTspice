* T2CU SPICE BSIM3 VERSION 3.1 PARAMETERS

* SPICE 3f5 Level 8, Star-HSPICE Level 49,* UTMOST Level 8

* DATE: Feb 18/03
* LOT: T2CU                  WAF: 0001
* Temperature_parameters=Default
.MODEL tsmc18N NMOS (                                LEVEL   = 8
+VERSION = 3.1            TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 2.3549E17      VTH0    = 0.3669193
+K1      = 0.592797       K2      = 2.518108E-3    K3      = 1E-3
+K3B     = 4.7942179      W0      = 1E-7           NLX     = 1.745125E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 1.3683195      DVT1    = 0.4097438      DVT2    = 0.0552615
+U0      = 263.5112775    UA      = -1.363381E-9   UB      = 2.253823E-18
+UC      = 4.833037E-11   VSAT    = 1.017805E5     A0      = 1.9261289
+AGS     = 0.4192338      B0      = -1.069507E-8   B1      = -1E-7
+KETA    = -8.579587E-3   A1      = 2.789024E-4    A2      = 0.8916186
+RDSW    = 126.5291844    PRWG    = 0.4957859      PRWB    = -0.2
+WR      = 1              WINT    = 0              LINT    = 7.790316E-9
+XL      = -2E-8          XW      = -1E-8          DWG     = -1.224589E-8
+DWB     = 1.579145E-8    VOFF    = -0.0895222     NFACTOR = 2.5
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 2.95614E-3     ETAB    = 1.374596E-4
+DSUB    = 0.013974       PCLM    = 0.7291486      PDIBLC1 = 0.1332365
+PDIBLC2 = 2.151668E-3    PDIBLCB = -0.1           DROUT   = 0.6947618
+PSCBE1  = 7.412661E10    PSCBE2  = 1.812826E-7    PVAG    = 9.540595E-3
+DELTA   = 0.01           RSH     = 5.9            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 8.71E-10       CGSO    = 8.71E-10       CGBO    = 1E-12
+CJ      = 9.67972E-4     PB      = 0.6966474      MJ      = 0.3609772
+CJSW    = 2.443898E-10   PBSW    = 0.8082076      MJSW    = 0.1013742
+CJSWG   = 3.3E-10        PBSWG   = 0.8082076      MJSWG   = 0.1013742
+CF      = 0              PVTH0   = 7.226579E-4    PRDSW   = -4.5298309
+PK2     = -4.696208E-4   WKETA   = 6.028223E-3    LKETA   = -8.791311E-3
+PU0     = 17.2549887     PUA     = 6.802365E-11   PUB     = 4.224871E-24
+PVSAT   = 1.298468E3     PETA0   = 1.003159E-4    PKETA   = -3.864603E-4    )
*
.MODEL tsmc18P PMOS (                                LEVEL   = 8 
+VERSION = 3.1            TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 4.1589E17      VTH0    = -0.4002789
+K1      = 0.5772615      K2      = 0.026742       K3      = 0
+K3B     = 14.2532769     W0      = 1E-6           NLX     = 9.883899E-8
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.6718731      DVT1    = 0.3118588      DVT2    = 0.1
+U0      = 118.0541064    UA      = 1.626518E-9    UB      = 1.229265E-21
+UC      = -1E-10         VSAT    = 2E5            A0      = 1.8109799
+AGS     = 0.4096261      B0      = 7.705744E-7    B1      = 2.657048E-6
+KETA    = 0.0212376      A1      = 0.5260122      A2      = 0.3207082
+RDSW    = 306.4304418    PRWG    = 0.5            PRWB    = 0.0612789
+WR      = 1              WINT    = 0              LINT    = 2.043723E-8
+XL      = -2E-8          XW      = -1E-8          DWG     = -4.602158E-8
+DWB     = 8.005928E-9    VOFF    = -0.0992452     NFACTOR = 2
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0.0331989      ETAB    = -0.0375363
+DSUB    = 0.7172358      PCLM    = 1.5224082      PDIBLC1 = 2.700462E-4
+PDIBLC2 = 0.0165863      PDIBLCB = -1E-3          DROUT   = 1.640424E-4
+PSCBE1  = 7.71553E9      PSCBE2  = 2.228426E-9    PVAG    = 5.1166248
+DELTA   = 0.01           RSH     = 6.7            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 6.92E-10       CGSO    = 6.92E-10       CGBO    = 1E-12
+CJ      = 1.173089E-3    PB      = 0.8524959      MJ      = 0.415401
+CJSW    = 2.217367E-10   PBSW    = 0.5936755      MJSW    = 0.2603391
+CJSWG   = 4.22E-10       PBSWG   = 0.5936755      MJSWG   = 0.2603391
+CF      = 0              PVTH0   = 1.425828E-3    PRDSW   = 0.9887283
+PK2     = 1.495689E-3    WKETA   = 0.0286138      LKETA   = -2.746502E-3
+PU0     = -1.2891258     PUA     = -5.395E-11     PUB     = 1E-21
+PVSAT   = -50            PETA0   = 1.003159E-4    PKETA   = -2.891811E-3    )
*
