.SUBCKT irl3714z_s_l 1 2 3
* Model generated on Jun 22, 04
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=2.63853 LAMBDA=0 KP=45.4893
+CGSO=4.45235e-06 CGDO=1.1492e-07
RS 8 3 0.0103197
D1 3 1 MD
.MODEL MD D IS=2.70143e-12 RS=0.00721606 N=1.04861 BV=20
+IBV=0.00025 EG=1.2 XTI=2.96785 TT=1.00001e-07
+CJO=2.76532e-10 VJ=0.5 M=0.409124 FC=0.5
RDS 3 1 1e+06
RD 9 1 0.0001
RG 2 7 2.18034
D2 4 5 MD1
.MODEL MD1 D IS=1e-32 N=50
+CJO=1.2665e-10 VJ=4.66779 M=0.3 FC=1e-08
D3 0 5 MD2
.MODEL MD2 D IS=1e-10 N=0.439082 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 4.35626e-10
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
.MODEL MD3 D IS=1e-10 N=0.439082
.ENDS irl3714z_s_l

*SPICE Thermal Model Subcircuit
.SUBCKT irl3714z_s_lt 3 0

R_RTHERM1         3 2  1.291698867 
R_RTHERM2         2 1  2.336748834
R_RTHERM3         1 0  0.651552298
C_CTHERM1         3 0  0.000104514
C_CTHERM2         2 0  0.000377447
C_CTHERM3         1 0  0.008398405

.ENDS irl3714z_s_lt 


