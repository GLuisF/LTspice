.SUBCKT irf7338 1 2 3 4 6 8
* DUAL N AND P CHANNEL MOSFET
* External Node Designations
* Node 1 -> N-channel Source
* Node 2 -> N-Channel Gate
* Node 3 -> P-Channel Source
* Node 4 -> P-Channel Gate
* Node 6 -> P-Channel Drain
* Node 8 -> N-Channel Drain
X1 8 2 1 irf7338-n
X2 6 4 3 irf7338-p
.ENDS irf7338

.SUBCKT irf7338-n 1 2 3
* SPICE3 MODEL WITH THERMAL RC NETWORK
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on May  6, 04
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=1.62693 LAMBDA=0.283092 KP=27.4025
+CGSO=4.71445e-06 CGDO=1e-11
RS 8 3 0.017538
D1 3 1 MD
.MODEL MD D IS=4.70825e-09 RS=0.0159221 N=1.5 BV=12
+IBV=0.00025 EG=1 XTI=1 TT=1e-07
+CJO=7.14086e-10 VJ=0.5 M=0.400706 FC=0.5
RDS 3 1 1e+06
RD 9 1 0.0001
RG 2 7 10.7454
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=3.32678e-10 VJ=1.54419 M=0.550127 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.417155 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 4.92353e-10
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.417155
.ENDS irf7338-n

*SPICE Thermal Model Subcircuit
.SUBCKT irf7338-nt 3 0

R_RTHERM1         3 2  5.943519682
R_RTHERM2         2 1  31.91794773
R_RTHERM3         1 0  24.64185115
C_CTHERM1         3 0  0.000224278
C_CTHERM2         2 0  0.014225852
C_CTHERM3         1 0  0.372131133

.ENDS irf7338-nt

.SUBCKT irf7338-p 1 2 3
* SPICE3 MODEL WITH THERMAL RC NETWORK
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on May  6, 04
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM PMOS LEVEL=1 IS=1e-32
+VTO=-1 LAMBDA=0.00128145 KP=14.1121
+CGSO=4.42693e-06 CGDO=1.54773e-08
RS 8 3 0.0001
D1 1 3 MD
.MODEL MD D IS=3.40041e-08 RS=0.0752214 N=1.5 BV=12
+IBV=0.00025 EG=1 XTI=3.08416 TT=1e-07
+CJO=2.09433e-10 VJ=0.5 M=0.687905 FC=0.307532
RDS 3 1 1e+06
RD 9 1 0.0614104
RG 2 7 40.6993
D2 5 4 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=2.36837e-10 VJ=0.5 M=0.393836 FC=1e-08
D3 5 0 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.4 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 2.36837e-10
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 6 0 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.4
.ENDS irf7338-p

*SPICE Thermal Model Subcircuit
.SUBCKT irf7338-pt 3 0

R_RTHERM1         3 2  7.835568501
R_RTHERM2         2 1  28.08073974
R_RTHERM3         1 0  26.57859385
C_CTHERM1         3 0  0.000128517
C_CTHERM2         2 0  0.014108247
C_CTHERM3         1 0  0.278419545

.ENDS irf7338-pt



