* AD811 SPICE Macro-model                   7/91, Rev. A   
*                                           JCB / PMI
*
*
* Copyright 1991 by Analog Devices, Inc.
*
* Refer to "README.DOC" file for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*              non-inverting input
*              | inverting input
*              | | positive supply
*              | | |  negative supply
*              | | |  |  output
*              | | |  |  |
.SUBCKT AD811  1 2 99 50 28
*
* INPUT STAGE
*
R1   99  8     1E3
R2   10 50     1E3
V1   99  9     11
D1   9   8     DX
V2   11 50     11
D2   10 11     DX
I1   99  5     920E-6
I2   4  50     920E-6
Q1   5   5  3  QN
Q2   4   4  3  QP
Q3   8   5 30  QN
Q4   10  4 30  QP
*
* INPUT ERROR SOURCES
* 
GB1  99  1     POLY(1)  1  22  2E-6  1E-6
GB2  99 30     POLY(1)  1  22  2E-6  1E-6
VOS  3   1     500E-6
LS1  30  2     4E-8
CS1  99  2     0.5E-12
CS2  50  2     0.5E-12
CIN  1  50     2E-12
*
EREF 97  0     22  0  1
*
* GAIN STAGE & DOMINANT POLE
*
R5   12 97     1.5E6
C3   12 97     3.9E-12
G1   97 12     99  8  1E-3
G2   12 97     10 50  1E-3
V3   99 13     2.9
V4   14 50     2.9
D3   12 13     DX
D4   14 12     DX
*
* POLE AT 400 MHZ
*
R8  17 97     1E6
C4  17 97     0.530E-15
G4  97 17     12 22  1E-6
*
* ZERO AT 150 MHZ
*
R20 18 19     1E6
R21 19 97     1
C20 18 19     -.530E-15
E20 18 97     17 22  1E6
*
* POLE AT 200 MHZ
*
R12 21 97     1E6
C8  21 97     0.395E-15
G8  97 21     19 22  1E-6
*
* OUTPUT STAGE
*
ISY 99 50     14.7E-3
R13 22 99     16.7E3
R14 22 50     16.7E3
R15 27 99     22
R16 27 50     22
L2  27 28     1E-8
G9  25 50     21 27  45.45E-3
G10 26 50     27 21  45.45E-3
G11 27 99     99 21  45.45E-3
G12 50 27     21 50  45.45E-3
V5  23 27     1.3
V6  27 24     1.3
D5  21 23     DX
D6  24 21     DX
D7  99 25     DX
D8  99 26     DX
D9  50 25     DY
D10 50 26     DY
*
* MODELS USED
*
.MODEL QN   NPN(BF=1E9 IS=1E-15)
.MODEL QP   PNP(BF=1E9 IS=1E-15)
.MODEL DX   D(IS=1E-15)
.MODEL DY   D(IS=1E-15 BV=50)
.ENDS AD811
