*
.SUBCKT CD4043 VCC R S Q E GND

XU3         7 VCC R VCC GND GATE_2INPUT_HC_2I_NAND_PP_ST_0
XU2         8 VCC S VCC GND GATE_2INPUT_HC_2I_NAND_PP_ST_0
XU1         9 10 7 VCC GND GATE_2INPUT_HC_2I_NAND_PP_ST_1
XU13        10 8 9 VCC GND GATE_2INPUT_HC_2I_NAND_PP_ST_0
XU8         Q 10 E VCC GND BUFFER_0

.ENDS
********************************************************************************
*                                 NAND_FLIPFLOP
********************************************************************************

.SUBCKT GATE_2INPUT_HC_2I_NAND_PP_ST_0  Y A B VCC AGND
XU1 Y A B VCC AGND LOGIC_GATE_2PIN_OD_HC_2I_NAND_PP_ST
.ENDS


*$
.SUBCKT LOGIC_GATE_2PIN_OD_HC_2I_NAND_PP_ST OUT A B VCC GND
.PARAM VCC_ABS_MAX = 20
.PARAM VCC_MAX = 6
.PARAM RA = 240000000
.PARAM RB = 240000000
.PARAM CA = 5E-15
.PARAM CB = 5E-15
.PARAM ROEZ = 5000
.PARAM COEZ = 3E-12
RA  A  GND {RA}
RB  B  GND {RB}
CA  A  GND {CA}
CB  B  GND {CB}
XUA NA A VCC GND LOGIC_INPUT_HC_2I_NAND_PP_ST
XUB NB B VCC GND LOGIC_INPUT_HC_2I_NAND_PP_ST
XUG NA NB NOUTG VCC GND LOGIC_FUNCTION_2_HC_2I_NAND_PP_ST
XUOUT NOUTG NOUT_INT VCC GND LOGIC_PP_OUTPUT_HC_2I_NAND_PP_ST
XICC VCC GND NVIOUT LOGIC_ICC_HC_2I_NAND_PP_ST
SICC VCC GND VCC GND SW1
* MONITOR OUTPUT CURRENT *
H1 NVIOUT GND VIOUT 1
VIOUT NOUT_INT OUTSW 0
SIOFF OUTSW OUT VCC GND SW2
.MODEL SW1 VSWITCH VON = {VCC_ABS_MAX} VOFF = {VCC_MAX} RON = 10 ROFF = 60E6
.MODEL SW2 VSWITCH VON = {0.55} VOFF = {0.45} RON = 10M ROFF = 100E6
.ENDS
*$

.SUBCKT LOGIC_INPUT_HC_2I_NAND_PP_ST OUT IN VCC VEE
ESTD_THR VSTD_THR VEE TABLE {V(VCC,VEE)} =
+(1,0.5)
+(6,3)
** OUTPUT VOLTAGES **
***********************************
**** STANDARD INPUT MODEL *********
***********************************
GSTD VEE CURR_OUT VALUE = {0.5*V(VCC,VEE)*(SGN(V(IN,VSTD_THR)) + ABS(SGN(V(IN,VSTD_THR))))}
ROUT CURR_OUT VEE 1
EMID MID VEE VALUE = {0.5*(V(VCC,VEE) + V(VEE))}
EARG NARG VEE VALUE = {V(CURR_OUT,VEE) - V(MID,VEE)}
EOUT OUT VEE VALUE = {0.5*(SGN(V(NARG,VEE)) + ABS(SGN(V(NARG,VEE) ) ) )}
*EOUT OUT VEE CURR_OUT VEE 1
.ENDS


*$
.SUBCKT LOGIC_FUNCTION_2_HC_2I_NAND_PP_ST A B OUT VCC VEE
GNAND VEE N1 VALUE = {(1 - V(A,VEE)*V(B,VEE))}
RN1 N1 VEE 1
EOUT OUT VEE N1 VEE 1
.ENDS


*$
.SUBCKT LOGIC_PP_OUTPUT_HC_2I_NAND_PP_ST IN OUT VCC VEE
EROH NROH VEE TABLE {V(VCC,VEE)} =
+(2,1)
+(6,1)
EROL NROL VEE TABLE {V(VCC,VEE)} =
+(2,1)
+(6,1)
E1 N1 VEE VALUE = {V(VCC,VEE)*V(IN,VEE)}
GOUT N1 OUT VALUE = {V(N1,OUT)*(V(IN,VEE)/V(NROH,VEE) + (1 - V(IN,VEE))/V(NROL,VEE))}
.ENDS
*


.SUBCKT LOGIC_ICC_HC_2I_NAND_PP_ST VCC VEE VIOUT
.PARAM ICC = 2.5E-08
.PARAM VCC_MAX = 6
.PARAM VCC_MIN = 2
*GICC VCC VEE VALUE = {ICC*V(VCC,VEE)/VCC_MAX}
GICC VCC VEE VALUE = {ICC*0.5*(1 + SGN(V(VCC,VEE) - VCC_MIN))}
*
* FLOATING GROUND AT MID-RAIL
EGNDF GNDF 0 VALUE = {0.5*(V(VCC) + V(VEE))}
*
GOUTP VCC GNDF VALUE = {V(VIOUT,VEE)*0.5*(SGN(V(VIOUT,VEE)) + ABS(SGN(V(VIOUT,VEE))))}
GOUTN GNDF VEE VALUE = {V(VIOUT,VEE)*0.5*(SGN(V(VIOUT,VEE)) + ABS(SGN(V(VIOUT,VEE))))}
*
*GOUTP VCC GNDF VALUE = {IF(V(VIMON,GNDF) > 0, V(VIMON,GNDF),0)}
*GOUTN GNDF VEE VALUE = {IF(V(VIMON,GNDF) <= 0, V(VIMON,GNDF),0)}
.ENDS
*$


********************************************************************************
*                                 NAND_FLIPFLOP
********************************************************************************

.SUBCKT GATE_2INPUT_HC_2I_NAND_PP_ST_1  Y A B VCC AGND
XU1 Y A B VCC AGND LOGIC_GATE_2PIN_OD_HC_2I_NAND_PP_ST_1
.ENDS


*$
.SUBCKT LOGIC_GATE_2PIN_OD_HC_2I_NAND_PP_ST_1 OUT A B VCC GND
.PARAM VCC_ABS_MAX = 20
.PARAM VCC_MAX = 6
.PARAM RA = 240000000
.PARAM RB = 240000000
.PARAM CA = 5E-15
.PARAM CB = 5E-15
.PARAM ROEZ = 5000
.PARAM COEZ = 3E-12
RA  A  GND {RA}
RB  B  GND {RB}
CA  A  GND {CA}
CB  B  GND {CB}
XUA NA A VCC GND LOGIC_INPUT_HC_2I_NAND_PP_ST
XUB NB B VCC GND LOGIC_INPUT_HC_2I_NAND_PP_ST
XUG NA NB NOUTG VCC GND LOGIC_FUNCTION_2_HC_2I_NAND_PP_ST
XUOUT NOUTG NOUT_INT VCC GND LOGIC_PP_OUTPUT_HC_2I_NAND_PP_ST_1
XICC VCC GND NVIOUT LOGIC_ICC_HC_2I_NAND_PP_ST
SICC VCC GND VCC GND SW1
* MONITOR OUTPUT CURRENT *
H1 NVIOUT GND VIOUT 1
VIOUT NOUT_INT OUTSW 0
SIOFF OUTSW OUT VCC GND SW2
.MODEL SW1 VSWITCH VON = {VCC_ABS_MAX} VOFF = {VCC_MAX} RON = 10 ROFF = 60E6
.MODEL SW2 VSWITCH VON = {0.55} VOFF = {0.45} RON = 10M ROFF = 100E6
.ENDS
*$


*$
.SUBCKT LOGIC_PP_OUTPUT_HC_2I_NAND_PP_ST_1 IN OUT VCC VEE
EROH NROH VEE TABLE {V(VCC,VEE)} =
+(2,10)
+(6,10)
EROL NROL VEE TABLE {V(VCC,VEE)} =
+(2,10)
+(6,10)
E1 N1 VEE VALUE = {V(VCC,VEE)*V(IN,VEE)}
GOUT N1 OUT VALUE = {V(N1,OUT)*(V(IN,VEE)/V(NROH,VEE) + (1 - V(IN,VEE))/V(NROL,VEE))}
.ENDS
*


********************************************************************************
*                                 TRI-STATE BUFFER
********************************************************************************

.SUBCKT BUFFER_0  Y A OEZ VCC AGND
XU1 Y A VCC OEZ VCC AGND LOGIC_GATE_2PIN_TRI_STATE_HC_1I_AND_TRISTATE_CMOS
.ENDS




.SUBCKT LOGIC_GATE_2PIN_TRI_STATE_HC_1I_AND_TRISTATE_CMOS OUT A B OEZ VCC GND
.PARAM VCC_ABS_MAX = 20
.PARAM VCC_MAX = 5.5
.PARAM RA = 220000000
.PARAM CA = 1E-11
.PARAM ROEZ = 5000
.PARAM COEZ = 3E-12
RA  A  GND {RA}
CA  A  GND {CA}
ROEZ OEZ GND {ROEZ}
COEZ OEZ GND {COEZ}
XUA NA A VCC GND LOGIC_INPUT_HC_1I_AND_TRISTATE_CMOS
XUB NB B VCC GND LOGIC_INPUT_HC_1I_AND_TRISTATE_CMOS
XUOEZ NOEZ OEZ VCC GND LOGIC_INPUT_HC_1I_AND_TRISTATE_CMOS
XUG NA NB NOUTG VCC GND LOGIC_FUNCTION_2_HC_1I_AND_TRISTATE_CMOS
XOUTPD NOUTG NOUTTPD VCC GND TPD_LVC_1i_AND_Tristate_CMOS
XUOUT NOUTTPD NOUT_INT NOEZ VCC GND LOGIC_TRI_STATE_OUTPUT_HC_1I_AND_TRISTATE_CMOS
XICC VCC GND NVIOUT LOGIC_ICC_HC_1I_AND_TRISTATE_CMOS
SICC VCC GND VCC GND SW1
H1 NVIOUT GND VIOUT 1
VIOUT NOUT_INT OUTSW 0
SIOFF OUTSW OUT VCC GND SW2
DA2 GND A D1
DB2 GND B D1
DO2 GND OUT D1
DOE1 NOEZ VCC D1
DOE2 GND OEZ D1
RDA1 NA1 GND 1E6
RDB1 NB1 GND 1E6
RDO1 NO1 GND 1E6
.MODEL SW1 VSWITCH VON = {VCC_ABS_MAX} VOFF = {VCC_MAX} RON = 10 ROFF = 60E6
.MODEL SW2 VSWITCH VON = {0.55} VOFF = {0.45} RON = 10M ROFF = 100E6
.MODEL D1 D
.ENDS


.SUBCKT LOGIC_INPUT_HC_1I_AND_TRISTATE_CMOS OUT IN VCC VEE
.PARAM STANDARD_INPUT_SELECT = 1
.PARAM SCHMITT_TRIGGER_INPUT_SELECT = 0
ESTD_THR VSTD_THR VEE TABLE {V(VCC,VEE)} =
+(1,0.5)
+(6,3)
GSTD VEE CURR_OUT VALUE = {STANDARD_INPUT_SELECT*0.5*V(VCC,VEE)*(SGN(V(IN,VSTD_THR)) + ABS(SGN(V(IN,VSTD_THR))))}
ROUT CURR_OUT VEE 1
EMID MID VEE VALUE = {0.5*(V(VCC,VEE) + V(VEE))}
EARG NARG VEE VALUE = {V(CURR_OUT,VEE) - V(MID,VEE)}
EOUT OUT VEE VALUE = {0.5*(SGN(V(NARG,VEE)) + ABS(SGN(V(NARG,VEE) ) ) )}
*EOUT OUT VEE CURR_OUT VEE 1
.ENDS

.SUBCKT LOGIC_FUNCTION_2_HC_1I_AND_TRISTATE_CMOS A B OUT VCC VEE
GAND  VEE N1 VALUE = {V(A,VEE)*V(B,VEE)}
RN1 N1 VEE 1
EOUT OUT VEE N1 VEE 1
.ENDS



.SUBCKT LOGIC_TRI_STATE_OUTPUT_HC_1I_AND_TRISTATE_CMOS IN OUT OEZ VCC VEE
EROH NROH VEE TABLE {V(VCC,VEE)} =
+(5,400)
+(10,192)
+(15,220)
EROL NROL VEE TABLE {V(VCC,VEE)} =
+(5,400)
+(10,192)
+(15,220)
EOEZ N2 VEE VALUE = {V(OEZ,VEE)}
E1 N1 VEE VALUE = {V(VCC,VEE)*V(IN,VEE)*V(N2,VEE)}
GOUT N1 OUT VALUE = {V(N1,OUT)*V(N2,VEE)*(V(IN,VEE)/V(NROH,VEE) + (1 - V(IN,VEE))/V(NROL,VEE))}
.ENDS

.SUBCKT  TPD_LVC_1i_AND_Tristate_CMOS IN OUT VCC VEE
.PARAM TPDELAY1 = 1N
.PARAM RS = 10K
.PARAM CS = {-TPDELAY1/(RS*LOG(0.5))}
*ETPDNORM NTPDNORM VEE TABLE {V(VCC,VEE)} =
*+({VCC1},{TPDELAY1/TPDELAY4})
*+({VCC2},{TPDELAY2/TPDELAY4})
*+({VCC3},{TPDELAY3/TPDELAY4})
*+({VCC4},{TPDELAY4/TPDELAY4})
ETPDNORM NTPDNORM VEE TABLE {V(VCC,VEE)} =
+(5,80)
+(10,25)
+(15,10)
*R1 IN N1 {RS}
G1 IN N1 VALUE = {V(IN,N1)/(V(NTPDNORM,VEE)*RS)}
RZ IN N1 10G
C1 N1 VEE {CS}
E1 N2 VEE VALUE = {0.5*(1 + SGN(V(N1,VEE) - 0.5))}
EOUT OUT VEE N2 VEE 1
.ENDS

.SUBCKT LOGIC_ICC_HC_1I_AND_TRISTATE_CMOS VCC VEE VIOUT
.PARAM ICC = 2.5E-07
.PARAM VCC_MAX = 5.5
.PARAM VCC_MIN = 2
GICC VCC VEE VALUE = {ICC*0.5*(1 + SGN(V(VCC,VEE) - VCC_MIN))}
EGNDF GNDF 0 VALUE = {0.5*(V(VCC) + V(VEE))}
GOUTP VCC GNDF VALUE = {V(VIOUT,VEE)*0.5*(SGN(V(VIOUT,VEE)) + ABS(SGN(V(VIOUT,VEE))))}
GOUTN GNDF VEE VALUE = {V(VIOUT,VEE)*0.5*(SGN(V(VIOUT,VEE)) + ABS(SGN(V(VIOUT,VEE))))}
.ENDS
